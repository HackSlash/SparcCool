// First test package

module SparCool;

initial begin
	$display("Hello World!");
	#10 $finish;
end

endmodule